library ieee;
use ieee.std_logic_1164.all;

entity tbird_lights is

port (L, R, H, CLK: in std_logic;
		LC,LB,LA,RA,RB,RC: out std_logic
);

end entity;


architecture behavioral of tbird_lights is

type STATE_TYPE is (s0, s1,s2,s3,s4,s5,s6,s7);
signal CURRENT_STATE, NEXT_STATE : STATE_TYPE;



begin

process(CURRENT_STATE, L,R,H)
variable INPUTS : std_logic_vector(2 downto 0);

begin
INPUTS := L&R&H;

case CURRENT_STATE is
when S0 => if(INPUTS = "000") then
			NEXT_STATE <= S0;
			elsif (INPUTS ="100") then
			NEXT_STATE <= S1;
			elsif (INPUTS = "010") then
			NEXT_STATE <= S4;
			else
			NEXT_STATE <= S7;
			end if;
			
when S1 => if(INPUTS(0) = '1') then
			NEXT_STATE <= S7;
			elsif (INPUTS ="100") then
			NEXT_STATE <= S2;
			else
			NEXT_STATE <= S0;
			end if;

when S2 => if(INPUTS(0) = '1') then
			NEXT_STATE <= S7;
			elsif (INPUTS ="100") then
			NEXT_STATE <= S3;
			else
			NEXT_STATE <= S0;
			end if;


when S3|S6 => if(INPUTS(0) = '1') then
			NEXT_STATE <= S7;
			elsif (INPUTS ="010") then
			NEXT_STATE <= S5;
			else
			NEXT_STATE <= S0;
			end if;


when S4 => if(INPUTS(0) = '1') then
			NEXT_STATE <= S7;
			elsif (INPUTS ="010") then
			NEXT_STATE <= S5;
			else
			NEXT_STATE <= S0;
			end if;


when S5 => if(INPUTS(0) = '1') then
			NEXT_STATE <= S7;
			elsif (INPUTS ="010") then
			NEXT_STATE <= S6;
			else
			NEXT_STATE <= S0;
			end if;


when S7 => NEXT_STATE <= S0;

end case;
end process;

process(CLK)
begin
	if (CLK'event and CLK = '1') then
	CURRENT_STATE <= NEXT_STATE;
	end if;
end process;
process(CURRENT_STATE)
begin
LC <= '0'; LB <= '0'; LA <= '0';
RA <= '0'; RB <= '0'; RC <= '0';
case CURRENT_STATE is

when S0 => null;
when S1 => LA <= '1';
when S2 => LA <= '1'; LB <= '1'; 
when S3 => LA <= '1'; LB <= '1'; LC <= '1';
when S4 => RA <= '1';
when S5 => RA <= '1'; RB <= '1';
when S6 => RA <= '1'; RB <= '1'; RC <= '1';
when S7 => LA <= '1'; LB <= '1'; LC <= '1';
			  RA <= '1'; RB <= '1'; RC <= '1';

end case;
end process;



end architecture;