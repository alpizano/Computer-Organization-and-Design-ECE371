library ieee;
use ieee.std_logic_1164.all;

entity 4to1_mux is

port ( s1 : in std_logic;
       s0 : in std_logic;
		 D3 : in std_logic;
		 D2 : in std_logic;
		 D1 : in std_logic;
		 D0 : in std_logic;
		 y  : out std_logic
     );



end entity 4to1_mux;

architecture dataflow of 4to1_mux is


begin

end architecture dataflow;