library ieee;
use ieee.std_logic_1164.all;

entity rotator_4bit is
port(A: in std_logic;
	  B: out std_logic
);


end entity rotator_4bit;

architecture dataflow of rotator_4bit is


begin


end architecture dataflow;